`timescale 10ns/1ns
module FPGA_EXP3_fhr_tb();
	reg a,res,c;
	wire out,e;
	wire [3:0]st;
	always begin
		#0 res=1'b0;c=1'b1;
		#100 res=1'b1;
		#10 a=1'b0;#10 a=1'b0;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
		#10 a=1'b0;#10 a=1'b1;
	end
	FPGA_EXP3_fhr U1(a,res,c,out,e,st);
endmodule